library verilog;
use verilog.vl_types.all;
entity tb_Huffman_Machine is
end tb_Huffman_Machine;
