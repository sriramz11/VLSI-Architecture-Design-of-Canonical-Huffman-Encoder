library verilog;
use verilog.vl_types.all;
entity tb_Canonical_Huffman_Machine is
end tb_Canonical_Huffman_Machine;
